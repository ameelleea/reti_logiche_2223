//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "it"
//: property prefix = "_GG"
//: property title = "mINV.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w13;    //: /sn:0 {0}(480,702)(205,702)(205,1056){1}
//: {2}(207,1058)(371,1058){3}
//: {4}(203,1058)(158,1058){5}
//: {6}(156,1056)(156,738)(351,738){7}
//: {8}(154,1058)(-49,1058)(-49,994)(-55,994){9}
//: {10}(-57,992)(-57,889)(-31,889){11}
//: {12}(-57,996)(-57,997)(-162,997){13}
supply0 w22;    //: /sn:0 {0}(527,923)(527,906)(488,906){1}
reg w12;    //: /sn:0 {0}(-162,840)(-143,840)(-143,840)(-128,840){1}
reg [3:0] w32;    //: /sn:0 {0}(#:267,674)(267,778)(349,778)(349,780){1}
reg [3:0] w33;    //: /sn:0 {0}(#:484,648)(484,665)(454,665)(454,690)(384,690)(384,710){1}
reg [3:0] w14;    //: /sn:0 {0}(#:392,674)(392,680)(438,680)(438,741){1}
reg [3:0] w5;    //: /sn:0 {0}(#:605,648)(605,665)(513,665)(513,674){1}
wire w6;    //: /sn:0 {0}(339,805)(43,805){1}
//: {2}(41,803)(41,766)(428,766){3}
//: {4}(41,807)(41,878){5}
//: {6}(39,880)(26,880){7}
//: {8}(41,882)(41,933){9}
//: {10}(39,935)(21,935){11}
//: {12}(41,937)(41,969)(389,969){13}
wire [3:0] w7;    //: /sn:0 {0}(#:398,873)(#:398,866)(367,866)(367,842){1}
//: {2}(367,838)(#:367,824){3}
//: {4}(#:365,840)(349,840)(349,871)(310,871)(310,861){5}
wire [3:0] w25;    //: /sn:0 {0}(#:386,780)(#:386,752){1}
wire [3:0] w0;    //: /sn:0 {0}(#:404,1030)(404,1024){1}
//: {2}(404,1020)(404,994){3}
//: {4}(#:402,1022)(321,1022)(321,1015){5}
wire [7:0] w30;    //: /sn:0 {0}(#:514,1146)(514,1179)(427,1179)(427,1145){1}
wire [3:0] w29;    //: /sn:0 {0}(#:515,716)(515,739)(475,739)(#:475,741){1}
wire w18;    //: /sn:0 {0}(-81,860)(-46,860){1}
//: {2}(-42,860)(-31,860){3}
//: {4}(-44,858)(-44,781){5}
wire [3:0] w10;    //: /sn:0 {0}(#:456,810)(456,800){1}
//: {2}(#:458,798)(496,798)(496,871)(528,871)(528,861){3}
//: {4}(456,796)(#:456,785){5}
wire [3:0] w23;    //: /sn:0 {0}(#:447,1102)(447,1055)(444,1055)(444,1023){1}
//: {2}(#:446,1021)(504,1021)(504,1015){3}
//: {4}(444,1019)(#:444,994){5}
wire w21;    //: /sn:0 {0}(-21,936)(-100,936){1}
//: {2}(-104,936)(-145,936)(-145,869)(-128,869){3}
//: {4}(-102,938)(-102,955)(-185,955)(-185,945){5}
wire [3:0] w1;    //: /sn:0 {0}(#:421,952)(#:421,939){1}
wire [3:0] w27;    //: /sn:0 {0}(#:406,1072)(#:406,1102){1}
wire [3:0] w9;    //: /sn:0 {0}(#:459,853)(#:459,873){1}
wire w26;    //: /sn:0 {0}(359,903)(366,903){1}
//: enddecls

  REG4 g8 (.in(w5), .clk(w13), .out(w29));   //: @(481, 675) /sz:(65, 40) /sn:0 /p:[ Ti0>1 Li0>0 Bo0<0 ]
  //: LED g44 (w7) @(310,854) /sn:0 /w:[ 5 ] /type:3
  //: joint g4 (w7) @(367, 840) /w:[ -1 2 4 1 ]
  //: DIP B (w14) @(392,664) /w:[ 0 ] /st:3 /dn:1
  //: joint g3 (w10) @(456, 798) /w:[ 2 4 -1 1 ]
  mAND g26 (.a(w12), .b(w21), .out0(w18));   //: @(-127, 821) /sz:(45, 68) /sn:0 /p:[ Li0>1 Li1>3 Ro0<0 ]
  DEMUX4 g2 (.A(w1), .c(w6), .ou1(w0), .ou2(w23));   //: @(390, 953) /sz:(66, 40) /sn:0 /p:[ Ti0>0 Li0>13 Bo0<3 Bo1<5 ]
  MUX4 g1 (.A(w14), .B(w29), .C(w6), .out(w10));   //: @(429, 742) /sz:(66, 42) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>3 Bo0<5 ]
  FFDet g24 (.D(w18), .Clk(w13), .Y(w6));   //: @(-30, 847) /sz:(55, 53) /sn:0 /p:[ Li0>3 Li1>11 Ro0<7 ]
  //: LED g39 (w21) @(-185,938) /sn:0 /w:[ 5 ] /type:0
  //: DIP A (w32) @(267,664) /w:[ 0 ] /st:10 /dn:1
  mINV g25 (.w1(w6), .w2(w21));   //: @(-20, 911) /sz:(40, 48) /R:2 /sn:0 /p:[ Ri0>11 Lo0<0 ]
  //: joint g10 (w6) @(41, 805) /w:[ 1 2 -1 4 ]
  //: LED g49 (w23) @(504,1008) /sn:0 /w:[ 3 ] /type:3
  //: SWITCH Clock (w13) @(-179,997) /w:[ 13 ] /st:0 /dn:1
  REG4 g6 (.in(w33), .clk(w13), .out(w25));   //: @(352, 711) /sz:(65, 40) /sn:0 /p:[ Ti0>1 Li0>7 Bo0<1 ]
  //: GROUND g35 (w22) @(527,929) /sn:0 /w:[ 0 ]
  //: joint g7 (w23) @(444, 1021) /w:[ 2 4 -1 1 ]
  //: joint g9 (w6) @(41, 880) /w:[ -1 5 6 8 ]
  COMPL2 g33 (.N(w10), .O(w9));   //: @(430, 811) /sz:(54, 41) /sn:0 /p:[ Ti0>0 Bo0<0 ]
  //: LED g45 (w30) @(514,1139) /sn:0 /w:[ 0 ] /type:3
  //: LED g41 (w10) @(528,854) /sn:0 /w:[ 3 ] /type:3
  MUL4 g42 (.A(w27), .B(w23), .out(w30));   //: @(386, 1103) /sz:(82, 41) /sn:0 /p:[ Ti0>1 Ti1>0 Bo0<1 ]
  //: joint g40 (w21) @(-102, 936) /w:[ 1 -1 2 4 ]
  //: joint g12 (w13) @(-57, 994) /w:[ 9 10 -1 12 ]
  RCA4 g34 (.A(w7), .B(w9), .cin(w22), .cout(w26), .S(w1));   //: @(367, 874) /sz:(120, 64) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  //: SWITCH g28 (w12) @(-179,840) /sn:0 /w:[ 0 ] /st:0 /dn:1
  REG4 g14 (.in(w0), .clk(w13), .out(w27));   //: @(372, 1031) /sz:(65, 40) /sn:0 /p:[ Ti0>0 Li0>3 Bo0<0 ]
  //: joint g5 (w0) @(404, 1022) /w:[ -1 2 4 1 ]
  //: joint g11 (w6) @(41, 935) /w:[ -1 9 10 12 ]
  //: DIP C (w33) @(484,638) /w:[ 0 ] /st:3 /dn:1
  //: DIP D (w5) @(605,638) /w:[ 0 ] /st:1 /dn:1
  MUX4 g0 (.A(w32), .B(w25), .C(w6), .out(w7));   //: @(340, 781) /sz:(66, 42) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Bo0<3 ]
  //: joint g38 (w18) @(-44, 860) /w:[ 2 4 1 -1 ]
  //: joint g15 (w13) @(156, 1058) /w:[ 5 6 8 -1 ]
  //: LED g37 (w18) @(-44,774) /sn:0 /w:[ 5 ] /type:0
  //: LED g53 (w0) @(321,1008) /sn:0 /w:[ 5 ] /type:3
  //: joint g13 (w13) @(205, 1058) /w:[ 2 1 4 -1 ]

endmodule
//: /netlistEnd

//: /netlistBegin FFDls
module FFDls(Y, Clk, D);
//: interface  /sz:(46, 61) /bd:[ Li0>D(9/61) Li1>Clk(49/61) Ro0<Y(36/61) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input Clk;    //: /sn:0 {0}(289,238)(274,238)(274,208){1}
//: {2}(274,204)(274,168)(289,168){3}
//: {4}(272,206)(143,206){5}
input D;    //: /sn:0 {0}(193,268)(175,268)(175,141){1}
//: {2}(177,139)(289,139){3}
//: {4}(173,139)(148,139){5}
output Y;    //: /sn:0 {0}(541,180)(493,180){1}
//: {2}(489,180)(469,180){3}
//: {4}(491,182)(491,229)(416,229)(416,254)(426,254){5}
wire w7;    //: /sn:0 {0}(426,288)(351,288)(351,258)(336,258){1}
wire w4;    //: /sn:0 {0}(425,159)(336,159){1}
wire w0;    //: /sn:0 {0}(470,275)(480,275)(480,221)(410,221)(410,193)(425,193){1}
wire w1;    //: /sn:0 {0}(235,267)(289,267){1}
//: enddecls

  //: joint g4 (D) @(175, 139) /w:[ 2 -1 4 1 ]
  mNOR g8 (.A(Y), .B(w7), .out(w0));   //: @(427, 238) /sz:(42, 64) /sn:0 /p:[ Li0>5 Li1>0 Ro0<0 ]
  mAND g3 (.a(Clk), .b(w1), .out0(w7));   //: @(290, 219) /sz:(45, 68) /sn:0 /p:[ Li0>0 Li1>1 Ro0<1 ]
  mAND g2 (.a(D), .b(Clk), .out0(w4));   //: @(290, 120) /sz:(45, 68) /sn:0 /p:[ Li0>3 Li1>3 Ro0<1 ]
  mINV g1 (.w1(D), .w2(w1));   //: @(194, 244) /sz:(40, 48) /sn:0 /p:[ Li0>0 Ro0<0 ]
  //: joint g10 (Y) @(491, 180) /w:[ 1 -1 2 4 ]
  //: joint g6 (Clk) @(274, 206) /w:[ -1 2 4 1 ]
  mNOR g7 (.A(w4), .B(w0), .out(Y));   //: @(426, 143) /sz:(42, 64) /sn:0 /p:[ Li0>0 Li1>1 Ro0<3 ]
  //: OUT g9 (Y) @(538,180) /sn:0 /w:[ 0 ]
  //: IN g5 (Clk) @(141,206) /sn:0 /w:[ 5 ]
  //: IN g0 (D) @(146,139) /sn:0 /w:[ 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin COMPL2
module COMPL2(O, N);
//: interface  /sz:(54, 41) /bd:[ Ti0>N[3:0](26/54) Bo0<O[3:0](29/54) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
supply1 w0;    //: /sn:0 {0}(754,310)(754,337)(714,337){1}
output [3:0] O;    //: /sn:0 {0}(#:529,575)(552,575)(#:552,477){1}
input [3:0] N;    //: /sn:0 {0}(#:314,54)(389,54){1}
//: {2}(390,54)(485,54){3}
//: {4}(486,54)(579,54){5}
//: {6}(580,54)(681,54){7}
//: {8}(682,54)(#:756,54){9}
wire w16;    //: /sn:0 {0}(456,334)(422,334){1}
wire w6;    //: /sn:0 {0}(580,311)(580,243){1}
wire w7;    //: /sn:0 {0}(579,201)(579,50){1}
wire w4;    //: /sn:0 {0}(390,309)(390,243){1}
wire w3;    //: /sn:0 {0}(484,199)(484,57)(485,57)(485,50){1}
wire w20;    //: /sn:0 {0}(567,471)(567,460)(685,460)(685,363){1}
wire w19;    //: /sn:0 {0}(347,333)(362,333){1}
wire w12;    //: /sn:0 {0}(682,312)(682,241){1}
wire w10;    //: /sn:0 {0}(547,471)(547,431)(487,431)(487,361){1}
wire w1;    //: /sn:0 {0}(389,201)(389,50){1}
wire w8;    //: /sn:0 {0}(484,310)(484,264)(485,264)(485,241){1}
wire w17;    //: /sn:0 {0}(583,362)(583,448)(557,448)(557,471){1}
wire w14;    //: /sn:0 {0}(654,336)(612,336){1}
wire w15;    //: /sn:0 {0}(537,471)(537,456)(393,456)(393,360){1}
wire w5;    //: /sn:0 {0}(681,199)(681,50){1}
wire w9;    //: /sn:0 {0}(516,335)(552,335){1}
//: enddecls

  assign w7 = N[1]; //: TAP g8 @(579,52) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  mINV g4 (.w1(w5), .w2(w12));   //: @(657, 200) /sz:(48, 40) /R:3 /sn:0 /p:[ Ti0>0 Bo0<1 ]
  //: OUT g16 (O) @(532,575) /sn:0 /R:2 /w:[ 0 ]
  mINV g3 (.w1(w3), .w2(w8));   //: @(460, 200) /sz:(48, 40) /R:3 /sn:0 /p:[ Ti0>0 Bo0<1 ]
  HA g17 (.N(w12), .cin(w0), .cout(w14), .S(w20));   //: @(655, 313) /sz:(58, 49) /sn:0 /p:[ Ti0>0 Ri0>1 Lo0<0 Bo0<1 ]
  mINV g2 (.w1(w1), .w2(w4));   //: @(365, 202) /sz:(48, 40) /R:3 /sn:0 /p:[ Ti0>0 Bo0<1 ]
  HA g1 (.N(w6), .cin(w14), .cout(w9), .S(w17));   //: @(553, 312) /sz:(58, 49) /sn:0 /p:[ Ti0>0 Ri0>1 Lo0<1 Bo0<0 ]
  HA g10 (.N(w8), .cin(w9), .cout(w16), .S(w10));   //: @(457, 311) /sz:(58, 49) /sn:0 /p:[ Ti0>0 Ri0>0 Lo0<0 Bo0<1 ]
  assign w1 = N[3]; //: TAP g6 @(389,52) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  assign w5 = N[0]; //: TAP g9 @(681,52) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  assign w3 = N[2]; //: TAP g7 @(485,52) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: VDD g12 (w0) @(765,310) /sn:0 /w:[ 0 ]
  HA g11 (.N(w4), .cin(w16), .cout(w19), .S(w15));   //: @(363, 310) /sz:(58, 49) /sn:0 /p:[ Ti0>0 Ri0>1 Lo0<1 Bo0<1 ]
  mINV g5 (.w1(w7), .w2(w6));   //: @(555, 202) /sz:(48, 40) /R:3 /sn:0 /p:[ Ti0>0 Bo0<1 ]
  //: IN g0 (N) @(758,54) /sn:0 /R:2 /w:[ 9 ]
  assign O = {w15, w10, w17, w20}; //: CONCAT g13  @(552,476) /sn:0 /R:3 /w:[ 1 0 0 1 0 ] /dr:1 /tp:0 /drp:1

endmodule
//: /netlistEnd

//: /netlistBegin DEMUX
module DEMUX(ou2, ou1, c, A);
//: interface  /sz:(63, 40) /bd:[ Ti0>A(30/63) Li0>c(16/40) Bo0<ou2(52/63) Bo1<ou1(12/63) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input A;    //: /sn:0 {0}(349,334)(177,334)(177,230)(169,230){1}
//: {2}(167,228)(167,165)(345,165){3}
//: {4}(167,232)(167,234)(138,234){5}
output ou2;    //: /sn:0 {0}(396,325)(426,325)(426,308)(441,308){1}
output ou1;    //: /sn:0 {0}(392,185)(421,185)(421,230)(436,230){1}
input c;    //: /sn:0 {0}(138,308)(226,308){1}
//: {2}(230,308)(336,308)(336,305)(349,305){3}
//: {4}(228,306)(228,197)(241,197){5}
wire w0;    //: /sn:0 {0}(283,196)(327,196)(327,194)(345,194){1}
//: enddecls

  mAND g4 (.b(w0), .a(A), .out0(ou1));   //: @(346, 146) /sz:(45, 68) /sn:0 /p:[ Li0>1 Li1>3 Ro0<0 ]
  //: joint g8 (c) @(228, 308) /w:[ 2 4 1 -1 ]
  //: OUT g3 (ou2) @(438,308) /sn:0 /w:[ 1 ]
  //: OUT g2 (ou1) @(433,230) /sn:0 /w:[ 1 ]
  //: IN g1 (c) @(136,308) /sn:0 /w:[ 0 ]
  mINV g6 (.w1(c), .w2(w0));   //: @(242, 173) /sz:(40, 48) /sn:0 /p:[ Li0>5 Ro0<0 ]
  //: joint g7 (A) @(167, 230) /w:[ 1 2 -1 4 ]
  mAND g5 (.b(A), .a(c), .out0(ou2));   //: @(350, 286) /sz:(45, 68) /sn:0 /p:[ Li0>0 Li1>3 Ro0<0 ]
  //: IN g0 (A) @(136,234) /sn:0 /w:[ 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin mOR
module mOR(b, a, out);
//: interface  /sz:(42, 45) /bd:[ Li0>a(14/45) Li1>b(33/45) Ro0<out(27/45) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(50,264)(136,264)(136,237)(151,237){1}
output out;    //: /sn:0 {0}(345,223)(284,223){1}
input a;    //: /sn:0 {0}(44,177)(136,177)(136,203)(151,203){1}
wire w0;    //: /sn:0 {0}(195,224)(242,224){1}
//: enddecls

  //: IN g4 (b) @(48,264) /sn:0 /w:[ 0 ]
  //: IN g3 (a) @(42,177) /sn:0 /w:[ 0 ]
  mNOR g1 (.B(b), .A(a), .out(w0));   //: @(152, 187) /sz:(42, 64) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: OUT g5 (out) @(342,223) /sn:0 /w:[ 0 ]
  mINV g0 (.w1(w0), .w2(out));   //: @(243, 200) /sz:(40, 48) /sn:0 /p:[ Li0>1 Ro0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin REG4
module REG4(clk, out, in);
//: interface  /sz:(65, 40) /bd:[ Ti0>in[3:0](32/65) Li0>clk(27/40) Bo0<out[3:0](34/65) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [3:0] in;    //: /sn:0 {0}(#:79,127)(97,127)(97,147){1}
//: {2}(97,148)(97,231){3}
//: {4}(97,232)(97,338){5}
//: {6}(97,339)(97,438){7}
//: {8}(97,439)(97,473){9}
input clk;    //: /sn:0 {0}(79,512)(119,512)(119,470){1}
//: {2}(121,468)(144,468){3}
//: {4}(119,466)(119,370){5}
//: {6}(121,368)(144,368){7}
//: {8}(119,366)(119,263){9}
//: {10}(121,261)(144,261){11}
//: {12}(119,259)(119,177)(144,177){13}
output [3:0] out;    //: /sn:0 {0}(319,306)(#:273,306){1}
wire w6;    //: /sn:0 {0}(101,439)(122,439)(122,439)(144,439){1}
wire w4;    //: /sn:0 {0}(101,232)(122,232)(122,232)(144,232){1}
wire w1;    //: /sn:0 {0}(101,148)(144,148){1}
wire w8;    //: /sn:0 {0}(267,321)(252,321)(252,459)(201,459){1}
wire w2;    //: /sn:0 {0}(267,291)(253,291)(253,168)(201,168){1}
wire w11;    //: /sn:0 {0}(267,311)(216,311)(216,359)(201,359){1}
wire w5;    //: /sn:0 {0}(267,301)(216,301)(216,252)(201,252){1}
wire w9;    //: /sn:0 {0}(101,339)(122,339)(122,339)(144,339){1}
//: enddecls

  FFDet g4 (.D(w6), .Clk(clk), .Y(w8));   //: @(145, 426) /sz:(55, 53) /sn:0 /p:[ Li0>1 Li1>3 Ro0<1 ]
  assign w6 = in[3]; //: TAP g8 @(95,439) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  assign w1 = in[0]; //: TAP g3 @(95,148) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  FFDet g2 (.D(w4), .Clk(clk), .Y(w5));   //: @(145, 219) /sz:(55, 53) /sn:0 /p:[ Li0>1 Li1>11 Ro0<1 ]
  FFDet g1 (.D(w1), .Clk(clk), .Y(w2));   //: @(145, 135) /sz:(55, 53) /sn:0 /p:[ Li0>1 Li1>13 Ro0<1 ]
  //: joint g10 (clk) @(119, 468) /w:[ 2 4 -1 1 ]
  assign w4 = in[1]; //: TAP g6 @(95,232) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  assign w9 = in[2]; //: TAP g7 @(95,339) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  //: IN g9 (clk) @(77,512) /sn:0 /w:[ 0 ]
  //: joint g12 (clk) @(119, 261) /w:[ 10 12 -1 9 ]
  FFDet g5 (.D(w9), .Clk(clk), .Y(w11));   //: @(145, 326) /sz:(55, 53) /sn:0 /p:[ Li0>1 Li1>7 Ro0<1 ]
  //: joint g11 (clk) @(119, 368) /w:[ 6 8 -1 5 ]
  //: OUT g14 (out) @(316,306) /sn:0 /w:[ 0 ]
  //: IN g0 (in) @(77,127) /sn:0 /w:[ 0 ]
  assign out = {w8, w11, w5, w2}; //: CONCAT g13  @(272,306) /sn:0 /w:[ 1 0 0 0 0 ] /dr:1 /tp:0 /drp:1

endmodule
//: /netlistEnd

//: /netlistBegin HA
module HA(cin, S, cout, N);
//: interface  /sz:(58, 49) /bd:[ Ti0>N(27/58) Ri0>cin(24/49) Lo0<cout(23/49) Bo0<S(30/58) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input cin;    //: /sn:0 {0}(380,364)(315,364)(315,310){1}
//: {2}(315,306)(315,278)(381,278){3}
//: {4}(313,308)(300,308){5}
output cout;    //: /sn:0 {0}(500,355)(463,355)(463,355)(427,355){1}
output S;    //: /sn:0 {0}(500,269)(425,269){1}
input N;    //: /sn:0 {0}(380,335)(346,335)(346,253){1}
//: {2}(348,251)(381,251){3}
//: {4}(344,251)(300,251){5}
//: enddecls

  //: joint g4 (N) @(346, 251) /w:[ 2 -1 4 1 ]
  mAND g3 (.b(cin), .a(N), .out0(cout));   //: @(381, 316) /sz:(45, 68) /sn:0 /p:[ Li0>0 Li1>0 Ro0<1 ]
  mEXOR g2 (.a(N), .b(cin), .out(S));   //: @(382, 238) /sz:(42, 55) /sn:0 /p:[ Li0>3 Li1>3 Ro0<1 ]
  //: IN g1 (cin) @(298,308) /sn:0 /w:[ 5 ]
  //: OUT g6 (S) @(497,269) /sn:0 /w:[ 0 ]
  //: OUT g7 (cout) @(497,355) /sn:0 /w:[ 0 ]
  //: joint g5 (cin) @(315, 308) /w:[ -1 2 4 1 ]
  //: IN g0 (N) @(298,251) /sn:0 /w:[ 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin FFDet
module FFDet(Clk, Y, D);
//: interface  /sz:(55, 53) /bd:[ Li0>D(13/53) Li1>Clk(42/53) Ro0<Y(33/53) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input Clk;    //: /sn:0 {0}(94,307)(123,307){1}
//: {2}(127,307)(289,307)(289,228)(309,228){3}
//: {4}(125,305)(125,274){5}
input D;    //: /sn:0 {0}(94,161)(162,161){1}
output Y;    //: /sn:0 {0}(437,215)(357,215){1}
wire w0;    //: /sn:0 {0}(124,232)(124,201)(162,201){1}
wire w2;    //: /sn:0 {0}(210,188)(309,188){1}
//: enddecls

  mINV g4 (.w1(Clk), .w2(w0));   //: @(101, 233) /sz:(48, 40) /R:1 /sn:0 /p:[ Bi0>5 To0<0 ]
  FFDls g3 (.D(w2), .Clk(Clk), .Y(Y));   //: @(310, 179) /sz:(46, 61) /sn:0 /p:[ Li0>1 Li1>3 Ro0<1 ]
  FFDls g2 (.D(D), .Clk(w0), .Y(w2));   //: @(163, 152) /sz:(46, 61) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: IN g1 (Clk) @(92,307) /sn:0 /w:[ 0 ]
  //: OUT g6 (Y) @(434,215) /sn:0 /w:[ 0 ]
  //: joint g5 (Clk) @(125, 307) /w:[ 2 4 1 -1 ]
  //: IN g0 (D) @(92,161) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin RCA4
module RCA4(cin, S, B, A, cout);
//: interface  /sz:(120, 64) /bd:[ Ti0>A[3:0](31/120) Ti1>B[3:0](92/120) Ri0>cin(32/64) Lo0<cout(29/64) Bo0<S[3:0](54/120) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [3:0] B;    //: /sn:0 {0}(#:297,164)(360,164){1}
//: {2}(361,164)(457,164){3}
//: {4}(458,164)(540,164){5}
//: {6}(541,164)(644,164){7}
//: {8}(645,164)(708,164){9}
input [3:0] A;    //: /sn:0 {0}(#:297,121)(382,121){1}
//: {2}(383,121)(477,121){3}
//: {4}(478,121)(562,121){5}
//: {6}(563,121)(665,121){7}
//: {8}(666,121)(702,121){9}
input cin;    //: /sn:0 {0}(744,155)(754,155)(754,244)(682,244){1}
output cout;    //: /sn:0 {0}(348,248)(281,248)(281,303)(268,303)(268,315)(281,315){1}
output [3:0] S;    //: /sn:0 {0}(#:512,353)(512,410)(#:471,410){1}
wire w16;    //: /sn:0 {0}(645,168)(645,221){1}
wire w6;    //: /sn:0 {0}(458,168)(458,176)(457,176)(457,221){1}
wire w7;    //: /sn:0 {0}(478,125)(478,221){1}
wire w4;    //: /sn:0 {0}(376,274)(376,332)(497,332)(497,347){1}
wire w0;    //: /sn:0 {0}(442,248)(415,248)(415,244)(400,244){1}
wire w19;    //: /sn:0 {0}(658,274)(658,332)(527,332)(527,347){1}
wire w12;    //: /sn:0 {0}(563,125)(563,133)(564,133)(564,221){1}
wire w10;    //: /sn:0 {0}(630,248)(595,248)(595,244)(580,244){1}
wire w1;    //: /sn:0 {0}(361,168)(361,176)(363,176)(363,221){1}
wire w17;    //: /sn:0 {0}(666,125)(666,221){1}
wire w14;    //: /sn:0 {0}(556,274)(556,307)(517,307)(517,347){1}
wire w11;    //: /sn:0 {0}(541,168)(541,176)(543,176)(543,221){1}
wire w2;    //: /sn:0 {0}(383,125)(383,133)(384,133)(384,221){1}
wire w5;    //: /sn:0 {0}(528,248)(509,248)(509,244)(494,244){1}
wire w9;    //: /sn:0 {0}(470,274)(470,322)(507,322)(507,347){1}
//: enddecls

  assign w7 = A[2]; //: TAP g8 @(478,119) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: IN g4 (cin) @(742,155) /sn:0 /w:[ 0 ]
  assign S = {w4, w9, w14, w19}; //: CONCAT g16  @(512,352) /sn:0 /R:3 /w:[ 0 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  FA g3 (.a(w17), .b(w16), .cin(cin), .cout(w10), .S(w19));   //: @(631, 222) /sz:(50, 51) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: OUT g17 (S) @(474,410) /sn:0 /R:2 /w:[ 1 ]
  FA g2 (.a(w12), .b(w11), .cin(w10), .cout(w5), .S(w14));   //: @(529, 222) /sz:(50, 51) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FA g1 (.a(w7), .b(w6), .cin(w5), .cout(w0), .S(w9));   //: @(443, 222) /sz:(50, 51) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: IN g10 (B) @(295,164) /sn:0 /w:[ 0 ]
  assign w17 = A[0]; //: TAP g6 @(666,119) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  assign w2 = A[3]; //: TAP g9 @(383,119) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  assign w12 = A[1]; //: TAP g7 @(563,119) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  assign w11 = B[1]; //: TAP g12 @(541,162) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  assign w1 = B[3]; //: TAP g14 @(361,162) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  assign w16 = B[0]; //: TAP g11 @(645,162) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: IN g5 (A) @(295,121) /sn:0 /w:[ 0 ]
  FA g0 (.a(w2), .b(w1), .cin(w0), .cout(cout), .S(w4));   //: @(349, 222) /sz:(50, 51) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: OUT g15 (cout) @(278,315) /sn:0 /w:[ 1 ]
  assign w6 = B[2]; //: TAP g13 @(458,162) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin mNAND
module mNAND(out, b, a);
//: interface  /sz:(53, 64) /bd:[ Li0>a(14/64) Li1>b(49/64) Ro0<out(38/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(203,371)(282,371){1}
//: {2}(286,371)(303,371){3}
//: {4}(284,369)(284,211)(325,211){5}
supply0 w0;    //: /sn:0 {0}(311,456)(311,395)(317,395)(317,380){1}
output out;    //: /sn:0 {0}(317,290)(317,260){1}
//: {2}(319,258)(329,258)(329,257)(391,257){3}
//: {4}(317,256)(317,246)(311,246)(311,236){5}
//: {6}(313,234)(339,234)(339,220){7}
//: {8}(309,234)(278,234)(278,220){9}
supply1 w2;    //: /sn:0 {0}(278,203)(278,189)(309,189){1}
//: {2}(313,189)(339,189)(339,203){3}
//: {4}(311,187)(311,143){5}
input a;    //: /sn:0 {0}(203,298)(224,298){1}
//: {2}(228,298)(267,298)(267,298)(303,298){3}
//: {4}(226,296)(226,211)(264,211){5}
wire w4;    //: /sn:0 {0}(317,363)(317,335)(317,335)(317,307){1}
//: enddecls

  _GGNMOS #(2, 1) g4 (.Z(out), .S(w4), .G(a));   //: @(311,298) /sn:0 /w:[ 0 1 3 ]
  //: joint g8 (a) @(226, 298) /w:[ 2 4 1 -1 ]
  _GGPMOS #(2, 1) g3 (.Z(out), .S(w2), .G(a));   //: @(272,211) /sn:0 /w:[ 9 0 5 ]
  //: OUT g2 (out) @(388,257) /sn:0 /w:[ 3 ]
  //: IN g1 (b) @(201,371) /sn:0 /w:[ 0 ]
  //: GROUND g10 (w0) @(311,462) /sn:0 /w:[ 0 ]
  _GGNMOS #(2, 1) g6 (.Z(w4), .S(w0), .G(b));   //: @(311,371) /sn:0 /w:[ 0 1 3 ]
  //: joint g7 (w2) @(311, 189) /w:[ 2 4 1 -1 ]
  //: joint g9 (out) @(311, 234) /w:[ 6 -1 8 5 ]
  //: joint g12 (b) @(284, 371) /w:[ 2 4 1 -1 ]
  _GGPMOS #(2, 1) g5 (.Z(out), .S(w2), .G(b));   //: @(333,211) /sn:0 /w:[ 7 3 5 ]
  //: VDD g11 (w2) @(322,143) /sn:0 /w:[ 5 ]
  //: IN g0 (a) @(201,298) /sn:0 /w:[ 0 ]
  //: joint g13 (out) @(317, 258) /w:[ 2 4 -1 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin mAND
module mAND(out0, b, a);
//: interface  /sz:(45, 68) /bd:[ Li0>a(19/68) Li1>b(48/68) Ro0<out0(39/68) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(54,230)(82,230)(82,226)(97,226){1}
output out0;    //: /sn:0 {0}(328,200)(243,200){1}
input a;    //: /sn:0 {0}(54,170)(82,170)(82,191)(97,191){1}
wire w2;    //: /sn:0 {0}(201,201)(167,201)(167,215)(152,215){1}
//: enddecls

  //: OUT g4 (out0) @(325,200) /sn:0 /w:[ 0 ]
  mINV g3 (.w1(w2), .w2(out0));   //: @(202, 177) /sz:(40, 48) /sn:0 /p:[ Li0>0 Ro0<1 ]
  mNAND g2 (.a(a), .b(b), .out(w2));   //: @(98, 177) /sz:(53, 64) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 ]
  //: IN g1 (b) @(52,230) /sn:0 /w:[ 0 ]
  //: IN g0 (a) @(52,170) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin MUX
module MUX(out, C, B, A);
//: interface  /sz:(67, 40) /bd:[ Ti0>A(15/67) Ti1>B(47/67) Li0>C(19/40) Bo0<out(33/67) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(120,191)(216,191){1}
input A;    //: /sn:0 {0}(120,98)(215,98){1}
output out;    //: /sn:0 {0}(440,163)(369,163){1}
input C;    //: /sn:0 {0}(216,220)(121,220)(121,266)(134,266){1}
//: {2}(136,264)(136,262)(151,262){3}
//: {4}(136,268)(136,303)(120,303){5}
wire w1;    //: /sn:0 {0}(193,261)(194,261)(194,127)(215,127){1}
wire w2;    //: /sn:0 {0}(325,150)(277,150)(277,118)(262,118){1}
wire w5;    //: /sn:0 {0}(325,169)(278,169)(278,211)(263,211){1}
//: enddecls

  //: OUT g8 (out) @(437,163) /sn:0 /w:[ 0 ]
  mAND g4 (.b(C), .a(B), .out0(w5));   //: @(217, 172) /sz:(45, 68) /sn:0 /p:[ Li0>0 Li1>1 Ro0<1 ]
  mAND g3 (.b(w1), .a(A), .out0(w2));   //: @(216, 79) /sz:(45, 68) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 ]
  //: IN g2 (C) @(118,303) /sn:0 /w:[ 5 ]
  //: IN g1 (B) @(118,191) /sn:0 /w:[ 0 ]
  mOR g6 (.b(w5), .a(w2), .out(out));   //: @(326, 136) /sz:(42, 45) /sn:0 /p:[ Li0>0 Li1>0 Ro0<1 ]
  //: joint g7 (C) @(136, 266) /w:[ -1 2 1 4 ]
  mINV g5 (.w1(C), .w2(w1));   //: @(152, 238) /sz:(40, 48) /sn:0 /p:[ Li0>3 Ro0<0 ]
  //: IN g0 (A) @(118,98) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin MUX4
module MUX4(out, C, B, A);
//: interface  /sz:(66, 42) /bd:[ Ti0>A[3:0](9/66) Ti1>B[3:0](46/66) Li0>C(24/42) Bo0<out[3:0](27/66) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [3:0] B;    //: /sn:0 {0}(#:123,152)(282,152){1}
//: {2}(283,152)(393,152){3}
//: {4}(394,152)(493,152){5}
//: {6}(494,152)(604,152){7}
//: {8}(605,152)(697,152){9}
input [3:0] A;    //: /sn:0 {0}(#:121,111)(250,111){1}
//: {2}(251,111)(360,111){3}
//: {4}(361,111)(460,111){5}
//: {6}(461,111)(572,111){7}
//: {8}(573,111)(694,111){9}
output [3:0] out;    //: /sn:0 {0}(412,445)(395,445)(#:395,386){1}
input C;    //: /sn:0 {0}(116,249)(202,249){1}
//: {2}(204,247)(204,225)(235,225){3}
//: {4}(204,251)(204,309)(329,309){5}
//: {6}(333,309)(431,309){7}
//: {8}(435,309)(529,309)(529,225)(557,225){9}
//: {10}(433,307)(433,225)(446,225){11}
//: {12}(331,307)(331,225)(346,225){13}
wire w13;    //: /sn:0 {0}(605,156)(605,205){1}
wire w7;    //: /sn:0 {0}(390,380)(390,337)(400,337)(400,262)(380,262)(380,247){1}
wire w4;    //: /sn:0 {0}(394,156)(394,205){1}
wire w3;    //: /sn:0 {0}(380,380)(380,337)(269,337)(269,247){1}
wire w0;    //: /sn:0 {0}(283,156)(283,205){1}
wire w12;    //: /sn:0 {0}(573,115)(573,205){1}
wire w1;    //: /sn:0 {0}(251,115)(251,205){1}
wire w8;    //: /sn:0 {0}(461,115)(461,123)(462,123)(462,205){1}
wire w11;    //: /sn:0 {0}(400,380)(400,347)(480,347)(480,247){1}
wire w15;    //: /sn:0 {0}(410,380)(410,360)(591,360)(591,247){1}
wire w5;    //: /sn:0 {0}(361,115)(361,123)(362,123)(362,205){1}
wire w9;    //: /sn:0 {0}(494,156)(494,205){1}
//: enddecls

  MUX g8 (.A(w12), .B(w13), .C(C), .out(w15));   //: @(558, 206) /sz:(67, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>9 Bo0<1 ]
  MUX g4 (.A(w1), .B(w0), .C(C), .out(w3));   //: @(236, 206) /sz:(67, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>3 Bo0<1 ]
  //: joint g16 (C) @(204, 249) /w:[ -1 2 1 4 ]
  //: OUT g3 (out) @(409,445) /sn:0 /w:[ 0 ]
  //: joint g17 (C) @(433, 309) /w:[ 8 10 7 -1 ]
  //: IN g2 (C) @(114,249) /sn:0 /w:[ 0 ]
  //: IN g1 (B) @(121,152) /sn:0 /w:[ 0 ]
  //: joint g18 (C) @(331, 309) /w:[ 6 12 5 -1 ]
  assign w8 = A[2]; //: TAP g10 @(461,109) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  assign w1 = A[0]; //: TAP g6 @(251,109) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  assign w5 = A[1]; //: TAP g9 @(361,109) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  MUX g7 (.A(w8), .B(w9), .C(C), .out(w11));   //: @(447, 206) /sz:(67, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>11 Bo0<1 ]
  assign w13 = B[3]; //: TAP g12 @(605,150) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  assign w0 = B[0]; //: TAP g14 @(283,150) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  assign w12 = A[3]; //: TAP g11 @(573,109) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  MUX g5 (.A(w5), .B(w4), .C(C), .out(w7));   //: @(347, 206) /sz:(67, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>13 Bo0<1 ]
  assign out = {w15, w11, w7, w3}; //: CONCAT g19  @(395,385) /sn:0 /R:3 /w:[ 1 0 0 0 0 ] /dr:0 /tp:0 /drp:1
  assign w9 = B[2]; //: TAP g15 @(494,150) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: IN g0 (A) @(119,111) /sn:0 /w:[ 0 ]
  assign w4 = B[1]; //: TAP g13 @(394,150) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin mINV
module mINV(w1, w2);
//: interface  /sz:(40, 48) /bd:[ Li0>w1(24/48) Ro0<w2(23/48) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
supply1 w6;    //: /sn:0 {0}(629,171)(629,192)(646,192)(646,213){1}
supply0 w7;    //: /sn:0 {0}(640,341)(640,320)(646,320)(646,299){1}
input w1;    //: /sn:0 {0}(540,255)(615,255){1}
//: {2}(617,253)(617,221)(632,221){3}
//: {4}(617,257)(617,290)(632,290){5}
output w2;    //: /sn:0 {0}(646,230)(646,261){1}
//: {2}(648,263)(684,263){3}
//: {4}(646,265)(646,282){5}
//: enddecls

  //: IN g4 (w1) @(538,255) /sn:0 /w:[ 0 ]
  //: GROUND g3 (w7) @(640,347) /sn:0 /w:[ 0 ]
  //: VDD g2 (w6) @(640,171) /sn:0 /w:[ 0 ]
  _GGNMOS #(2, 1) g1 (.Z(w2), .S(w7), .G(w1));   //: @(640,290) /sn:0 /w:[ 5 1 5 ]
  //: OUT g6 (w2) @(681,263) /sn:0 /w:[ 3 ]
  //: joint g7 (w2) @(646, 263) /w:[ 2 1 -1 4 ]
  //: joint g5 (w1) @(617, 255) /w:[ -1 2 1 4 ]
  _GGPMOS #(2, 1) g0 (.Z(w2), .S(w6), .G(w1));   //: @(640,221) /sn:0 /w:[ 0 1 3 ]

endmodule
//: /netlistEnd

//: /netlistBegin MAC
module MAC(S, Aout, B, A, Sout, Cout, Bout, C);
//: interface  /sz:(68, 85) /bd:[ Ti0>A(55/68) Ti1>S(20/68) Ri0>B(26/85) Ri1>C(65/85) Lo0<Bout(18/85) Lo1<Cout(63/85) Bo0<Aout(15/68) Bo1<Sout(48/68) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(170,297)(159,297)(159,274)(165,274)(165,264)(172,264)(172,257){1}
//: {2}(174,255)(279,255){3}
//: {4}(170,255)(152,255){5}
//: {6}(148,255)(133,255){7}
//: {8}(150,257)(150,302)(170,302){9}
input A;    //: /sn:0 {0}(133,226)(183,226){1}
//: {2}(187,226)(279,226){3}
//: {4}(185,224)(185,169)(216,169){5}
//: {6}(185,228)(185,238)(200,238)(200,174)(216,174){7}
output Sout;    //: /sn:0 {0}(467,373)(423,373){1}
output Aout;    //: /sn:0 {0}(210,118)(200,118)(200,133)(252,133)(252,172)(237,172){1}
output Cout;    //: /sn:0 {0}(420,447)(397,447)(397,401){1}
output Bout;    //: /sn:0 {0}(244,334)(206,334)(206,300)(191,300){1}
input C;    //: /sn:0 {0}(379,294)(393,294)(393,349){1}
input S;    //: /sn:0 {0}(133,386)(250,386)(250,386)(370,386){1}
wire w2;    //: /sn:0 {0}(326,246)(355,246)(355,365)(370,365){1}
//: enddecls

  //: IN g4 (S) @(131,386) /sn:0 /w:[ 0 ]
  //: OUT g8 (Aout) @(207,118) /sn:0 /w:[ 0 ]
  //: IN g3 (B) @(131,255) /sn:0 /w:[ 7 ]
  //: IN g2 (A) @(131,226) /sn:0 /w:[ 0 ]
  FA g1 (.cin(C), .b(S), .a(w2), .cout(Cout), .S(Sout));   //: @(371, 350) /sz:(51, 50) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Bo0<1 Ro0<1 ]
  //: joint g10 (B) @(172, 255) /w:[ 2 -1 4 1 ]
  //: OUT g6 (Sout) @(464,373) /sn:0 /w:[ 0 ]
  //: OUT g7 (Cout) @(417,447) /sn:0 /w:[ 0 ]
  //: OUT g9 (Bout) @(241,334) /sn:0 /w:[ 0 ]
  _GGAND2 #(6) g12 (.I0(A), .I1(A), .Z(Aout));   //: @(227,172) /sn:0 /w:[ 5 7 1 ]
  //: IN g5 (C) @(377,294) /sn:0 /w:[ 0 ]
  //: joint g11 (A) @(185, 226) /w:[ 2 4 1 6 ]
  //: joint g14 (B) @(150, 255) /w:[ 5 -1 6 8 ]
  mAND g0 (.a(A), .b(B), .out0(w2));   //: @(280, 207) /sz:(45, 68) /sn:0 /p:[ Li0>3 Li1>3 Ro0<0 ]
  _GGAND2 #(6) g13 (.I0(B), .I1(B), .Z(Bout));   //: @(181,300) /sn:0 /w:[ 0 9 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin mNOR
module mNOR(B, out, A);
//: interface  /sz:(42, 64) /bd:[ Li0>A(16/64) Li1>B(50/64) Ro0<out(37/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
supply1 w6;    //: /sn:0 {0}(324,54)(324,97){1}
input B;    //: /sn:0 {0}(88,317)(155,317)(155,317)(221,317){1}
//: {2}(225,317)(357,317){3}
//: {4}(223,315)(223,195)(310,195){5}
supply0 w4;    //: /sn:0 {0}(329,361)(329,344){1}
//: {2}(331,342)(371,342)(371,326){3}
//: {4}(327,342)(295,342)(295,274){5}
input A;    //: /sn:0 {0}(88,105)(161,105)(161,105)(235,105){1}
//: {2}(239,105)(310,105){3}
//: {4}(237,107)(237,265)(281,265){5}
output out;    //: /sn:0 {0}(324,204)(324,216){1}
//: {2}(326,218)(447,218){3}
//: {4}(324,220)(324,240){5}
//: {6}(326,242)(371,242)(371,309){7}
//: {8}(322,242)(295,242)(295,257){9}
wire w0;    //: /sn:0 {0}(324,187)(324,114){1}
//: enddecls

  _GGNMOS #(2, 1) g4 (.Z(out), .S(w4), .G(A));   //: @(289,265) /sn:0 /w:[ 9 5 5 ]
  //: joint g8 (w4) @(329, 342) /w:[ 2 -1 4 1 ]
  _GGPMOS #(2, 1) g3 (.Z(out), .S(w0), .G(B));   //: @(318,195) /sn:0 /w:[ 0 0 5 ]
  _GGPMOS #(2, 1) g2 (.Z(w0), .S(w6), .G(A));   //: @(318,105) /sn:0 /w:[ 1 1 3 ]
  //: IN g1 (B) @(86,317) /sn:0 /w:[ 0 ]
  //: joint g10 (A) @(237, 105) /w:[ 2 -1 1 4 ]
  //: joint g6 (out) @(324, 242) /w:[ 6 5 8 -1 ]
  //: GROUND g7 (w4) @(329,367) /sn:0 /w:[ 0 ]
  //: VDD g9 (w6) @(335,54) /sn:0 /w:[ 0 ]
  //: OUT g12 (out) @(444,218) /sn:0 /w:[ 3 ]
  _GGNMOS #(2, 1) g5 (.Z(out), .S(w4), .G(B));   //: @(365,317) /sn:0 /w:[ 7 3 3 ]
  //: joint g11 (B) @(223, 317) /w:[ 2 4 1 -1 ]
  //: IN g0 (A) @(86,105) /sn:0 /w:[ 0 ]
  //: joint g13 (out) @(324, 218) /w:[ 2 1 -1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin mEXOR
module mEXOR(out, b, a);
//: interface  /sz:(42, 55) /bd:[ Li0>b(40/55) Li1>a(13/55) Ro0<out(31/55) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(245,276)(145,276)(145,394){1}
//: {2}(147,396)(155,396){3}
//: {4}(143,396)(130,396)(130,351)(122,351){5}
output out;    //: /sn:0 {0}(465,328)(384,328){1}
input a;    //: /sn:0 {0}(245,360)(137,360)(137,244){1}
//: {2}(139,242)(155,242){3}
//: {4}(137,240)(137,205)(122,205){5}
wire w7;    //: /sn:0 {0}(329,339)(315,339)(315,384)(300,384){1}
wire w4;    //: /sn:0 {0}(329,304)(315,304)(315,265)(300,265){1}
wire w0;    //: /sn:0 {0}(197,241)(245,241){1}
wire w1;    //: /sn:0 {0}(197,395)(245,395){1}
//: enddecls

  mINV g4 (.w1(b), .w2(w1));   //: @(156, 372) /sz:(40, 48) /sn:0 /p:[ Li0>3 Ro0<0 ]
  //: joint g8 (a) @(137, 242) /w:[ 2 4 -1 1 ]
  mINV g3 (.w1(a), .w2(w0));   //: @(156, 218) /sz:(40, 48) /sn:0 /p:[ Li0>3 Ro0<0 ]
  //: OUT g2 (out) @(462,328) /sn:0 /w:[ 0 ]
  //: IN g1 (b) @(120,351) /sn:0 /w:[ 5 ]
  mNAND g6 (.a(a), .b(w1), .out(w7));   //: @(246, 346) /sz:(53, 64) /sn:0 /p:[ Li0>0 Li1>1 Ro0<1 ]
  mNAND g7 (.a(w4), .b(w7), .out(out));   //: @(330, 290) /sz:(53, 64) /sn:0 /p:[ Li0>0 Li1>0 Ro0<1 ]
  //: joint g9 (b) @(145, 396) /w:[ 2 1 4 -1 ]
  mNAND g5 (.a(w0), .b(b), .out(w4));   //: @(246, 227) /sz:(53, 64) /sn:0 /p:[ Li0>1 Li1>0 Ro0<1 ]
  //: IN g0 (a) @(120,205) /sn:0 /w:[ 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin FA
module FA(cin, b, cout, S, a);
//: interface  /sz:(51, 50) /bd:[ Ti0>cin(22/51) Li0>b(36/50) Li1>a(15/50) Bo0<cout(26/51) Ro0<S(23/50) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(268,253)(278,253)(278,297)(216,297){1}
input cin;    //: /sn:0 {0}(268,129)(278,129)(278,176)(213,176){1}
output cout;    //: /sn:0 {0}(125,418)(95,418)(95,367){1}
input a;    //: /sn:0 {0}(121,100)(181,100)(181,151){1}
output S;    //: /sn:0 {0}(269,378)(187,378)(187,323){1}
wire w6;    //: /sn:0 {0}(108,323)(108,296)(156,296){1}
wire w3;    //: /sn:0 {0}(184,272)(184,202){1}
wire w2;    //: /sn:0 {0}(89,323)(89,175)(153,175){1}
//: enddecls

  HA g4 (.N(w3), .cin(b), .cout(w6), .S(S));   //: @(157, 273) /sz:(58, 49) /sn:0 /p:[ Ti0>0 Ri0>1 Lo0<1 Bo0<1 ]
  HA g3 (.N(a), .cin(cin), .cout(w2), .S(w3));   //: @(154, 152) /sz:(58, 49) /sn:0 /p:[ Ti0>1 Ri0>1 Lo0<1 Bo0<1 ]
  //: IN g2 (cin) @(266,129) /sn:0 /w:[ 0 ]
  //: IN g1 (b) @(266,253) /sn:0 /w:[ 0 ]
  mOR g6 (.a(w6), .b(w2), .out(cout));   //: @(78, 324) /sz:(45, 42) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  //: OUT g12 (cout) @(122,418) /sn:0 /w:[ 0 ]
  //: OUT g5 (S) @(266,378) /sn:0 /w:[ 0 ]
  //: IN g0 (a) @(119,100) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin DEMUX4
module DEMUX4(ou2, A, c, ou1);
//: interface  /sz:(66, 40) /bd:[ Ti0>A[3:0](31/66) Li0>c(16/40) Bo0<ou2[3:0](54/66) Bo1<ou1[3:0](14/66) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [3:0] A;    //: /sn:0 {0}(#:134,117)(188,117)(188,117)(249,117){1}
//: {2}(250,117)(376,117){3}
//: {4}(377,117)(497,117){5}
//: {6}(498,117)(623,117){7}
//: {8}(624,117)(690,117){9}
output [3:0] ou2;    //: /sn:0 {0}(475,469)(472,469)(472,469)(454,469)(#:454,408){1}
output [3:0] ou1;    //: /sn:0 {0}(323,469)(305,469)(#:305,408){1}
input c;    //: /sn:0 {0}(134,165)(194,165){1}
//: {2}(198,165)(325,165){3}
//: {4}(329,165)(448,165){5}
//: {6}(452,165)(580,165)(580,246)(593,246){7}
//: {8}(450,167)(450,246)(467,246){9}
//: {10}(327,167)(327,246)(346,246){11}
//: {12}(196,167)(196,246)(220,246){13}
wire w6;    //: /sn:0 {0}(449,402)(449,341)(399,341)(399,271){1}
wire w7;    //: /sn:0 {0}(300,402)(300,350)(359,350)(359,271){1}
wire w4;    //: /sn:0 {0}(377,121)(377,229){1}
wire w3;    //: /sn:0 {0}(290,402)(290,381)(233,381)(233,271){1}
wire w0;    //: /sn:0 {0}(250,121)(250,129)(251,129)(251,229){1}
wire w12;    //: /sn:0 {0}(498,121)(498,229){1}
wire w10;    //: /sn:0 {0}(320,402)(320,371)(606,371)(606,271){1}
wire w8;    //: /sn:0 {0}(624,121)(624,229){1}
wire w14;    //: /sn:0 {0}(310,402)(310,359)(480,359)(480,271){1}
wire w11;    //: /sn:0 {0}(469,402)(469,384)(646,384)(646,271){1}
wire w2;    //: /sn:0 {0}(439,402)(439,378)(273,378)(273,271){1}
wire w15;    //: /sn:0 {0}(459,402)(459,365)(520,365)(520,271){1}
//: enddecls

  assign w12 = A[1]; //: TAP g8 @(498,115) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  DEMUX g4 (.A(w12), .c(c), .ou1(w14), .ou2(w15));   //: @(468, 230) /sz:(63, 40) /sn:0 /p:[ Ti0>1 Li0>9 Bo0<1 Bo1<1 ]
  //: OUT g16 (ou2) @(472,469) /sn:0 /w:[ 0 ]
  DEMUX g3 (.A(w8), .c(c), .ou1(w10), .ou2(w11));   //: @(594, 230) /sz:(63, 40) /sn:0 /p:[ Ti0>1 Li0>7 Bo0<1 Bo1<1 ]
  //: IN g2 (A) @(132,117) /sn:0 /w:[ 0 ]
  DEMUX g1 (.A(w4), .c(c), .ou1(w7), .ou2(w6));   //: @(347, 230) /sz:(63, 40) /sn:0 /p:[ Ti0>1 Li0>11 Bo0<1 Bo1<1 ]
  //: joint g10 (c) @(450, 165) /w:[ 6 -1 5 8 ]
  assign w4 = A[2]; //: TAP g6 @(377,115) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: IN g9 (c) @(132,165) /sn:0 /w:[ 0 ]
  assign w0 = A[3]; //: TAP g7 @(250,115) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: joint g12 (c) @(196, 165) /w:[ 2 -1 1 12 ]
  assign ou2 = {w2, w6, w15, w11}; //: CONCAT g14  @(454,407) /sn:0 /R:3 /w:[ 1 0 0 0 0 ] /dr:1 /tp:0 /drp:1
  //: joint g11 (c) @(327, 165) /w:[ 4 -1 3 10 ]
  assign w8 = A[0]; //: TAP g5 @(624,115) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: OUT g15 (ou1) @(320,469) /sn:0 /w:[ 0 ]
  DEMUX g0 (.A(w0), .c(c), .ou1(w3), .ou2(w2));   //: @(221, 230) /sz:(63, 40) /sn:0 /p:[ Ti0>1 Li0>13 Bo0<1 Bo1<1 ]
  assign ou1 = {w3, w7, w14, w10}; //: CONCAT g13  @(305,407) /sn:0 /R:3 /w:[ 1 0 0 0 0 ] /dr:1 /tp:0 /drp:1

endmodule
//: /netlistEnd

//: /netlistBegin MUL4
module MUL4(B, A, out);
//: interface  /sz:(82, 41) /bd:[ Ti0>A[3:0](20/82) Ti1>B[3:0](61/82) Bo0<out[7:0](41/82) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [3:0] B;    //: /sn:0 {0}(#:-289,210)(-222,210){1}
//: {2}(-221,210)(-148,210){3}
//: {4}(-147,210)(-74,210){5}
//: {6}(-73,210)(-2,210){7}
//: {8}(-1,210)(72,210){9}
//: {10}(73,210)(145,210){11}
//: {12}(146,210)(219,210){13}
//: {14}(220,210)(292,210){15}
//: {16}(293,210)(365,210){17}
//: {18}(366,210)(440,210){19}
//: {20}(441,210)(513,210){21}
//: {22}(514,210)(585,210){23}
//: {24}(586,210)(656,210){25}
//: {26}(657,210)(729,210){27}
//: {28}(730,210)(802,210){29}
//: {30}(803,210)(876,210){31}
//: {32}(877,210)(#:892,210){33}
input [3:0] A;    //: /sn:0 {0}(#:902,176)(848,176){1}
//: {2}(847,176)(775,176){3}
//: {4}(774,176)(702,176){5}
//: {6}(701,176)(629,176){7}
//: {8}(628,176)(556,176){9}
//: {10}(555,176)(485,176){11}
//: {12}(484,176)(411,176){13}
//: {14}(410,176)(338,176){15}
//: {16}(337,176)(264,176){17}
//: {18}(263,176)(191,176){19}
//: {20}(190,176)(117,176){21}
//: {22}(116,176)(44,176){23}
//: {24}(43,176)(-29,176){25}
//: {26}(-30,176)(-102,176){27}
//: {28}(-103,176)(-176,176){29}
//: {30}(-177,176)(-249,176){31}
//: {32}(-250,176)(#:-289,176){33}
output [7:0] out;    //: /sn:0 {0}(301,689)(241,689)(#:241,668){1}
wire w16;    //: /sn:0 {0}(609,381)(609,353)(711,353)(711,339){1}
wire w13;    //: /sn:0 {0}(384,481)(384,419)(200,419)(200,339){1}
wire w7;    //: /sn:0 {0}(-82,529)(-82,349)(-240,349)(-240,339){1}
wire w58;    //: /sn:0 {0}(542,446)(542,431)(273,431)(273,339){1}
wire w65;    //: /sn:0 {0}(73,292)(73,214){1}
wire w34;    //: /sn:0 {0}(775,292)(775,180){1}
wire w50;    //: /sn:0 {0}(514,292)(514,214){1}
wire w59;    //: /sn:0 {0}(220,292)(220,214){1}
wire w39;    //: /sn:0 {0}(38,580)(38,634)(226,634)(226,662){1}
wire w62;    //: /sn:0 {0}(146,292)(146,214){1}
wire w72;    //: /sn:0 {0}(-102,292)(-102,180){1}
wire w56;    //: /sn:0 {0}(293,292)(293,214){1}
wire w22;    //: /sn:0 {0}(494,471)(521,471)(521,473)(527,473){1}
wire w82;    //: /sn:0 {0}(256,662)(256,633)(555,633)(555,499){1}
wire w20;    //: /sn:0 {0}(579,469)(601,469)(601,434){1}
wire w60;    //: /sn:0 {0}(191,292)(191,180){1}
wire w29;    //: /sn:0 {0}(442,475)(405,475)(405,481){1}
wire w30;    //: /sn:0 {0}(246,662)(246,629)(341,629)(341,577){1}
wire w71;    //: /sn:0 {0}(-73,292)(-73,214){1}
wire w42;    //: /sn:0 {0}(-79,580)(-79,639)(216,639)(216,662){1}
wire w37;    //: /sn:0 {0}(781,406)(784,406)(784,339){1}
wire w19;    //: /sn:0 {0}(573,408)(563,408)(563,446){1}
wire w12;    //: /sn:0 {0}(126,339)(126,353)(183,353)(183,478){1}
wire w66;    //: /sn:0 {0}(44,292)(44,180){1}
wire w10;    //: /sn:0 {0}(126,523)(126,392)(-93,392)(-93,339){1}
wire w63;    //: /sn:0 {0}(117,292)(117,180){1}
wire w84;    //: /sn:0 {0}(163,546)(196,546)(196,531){1}
wire w54;    //: /sn:0 {0}(338,292)(338,180){1}
wire w70;    //: /sn:0 {0}(328,524)(328,384)(-20,384)(-20,339){1}
wire w24;    //: /sn:0 {0}(-50,554)(10,554){1}
wire w21;    //: /sn:0 {0}(266,662)(266,639)(752,639)(752,432){1}
wire w31;    //: /sn:0 {0}(139,576)(139,629)(236,629)(236,662){1}
wire w32;    //: /sn:0 {0}(877,292)(877,215){1}
wire w68;    //: /sn:0 {0}(0,292)(0,222)(-1,222)(-1,214){1}
wire w53;    //: /sn:0 {0}(367,292)(367,222)(366,222)(366,214){1}
wire w8;    //: /sn:0 {0}(25,527)(25,441)(-167,441)(-167,339){1}
wire w46;    //: /sn:0 {0}(749,381)(749,366)(566,366)(566,339){1}
wire w52;    //: /sn:0 {0}(588,381)(588,348)(494,348)(494,339){1}
wire w17;    //: /sn:0 {0}(220,501)(275,501)(275,551)(313,551){1}
wire w27;    //: /sn:0 {0}(848,292)(848,180){1}
wire w44;    //: /sn:0 {0}(586,292)(586,214){1}
wire w75;    //: /sn:0 {0}(-176,292)(-176,180){1}
wire w80;    //: /sn:0 {0}(-110,553)(-134,553)(-134,645)(206,645)(206,662){1}
wire w33;    //: /sn:0 {0}(276,662)(276,645)(857,645)(857,339){1}
wire w35;    //: /sn:0 {0}(804,292)(804,222)(803,222)(803,214){1}
wire w67;    //: /sn:0 {0}(46,527)(46,353)(53,353)(53,339){1}
wire w49;    //: /sn:0 {0}(349,524)(349,508)(369,508){1}
wire w14;    //: /sn:0 {0}(457,448)(457,360)(421,360)(421,339){1}
wire w45;    //: /sn:0 {0}(557,292)(557,188)(556,188)(556,180){1}
wire w69;    //: /sn:0 {0}(-29,292)(-29,180){1}
wire w11;    //: /sn:0 {0}(629,292)(629,180){1}
wire w2;    //: /sn:0 {0}(702,292)(702,180){1}
wire w41;    //: /sn:0 {0}(658,292)(658,222)(657,222)(657,214){1}
wire w48;    //: /sn:0 {0}(412,292)(412,188)(411,188)(411,180){1}
wire w74;    //: /sn:0 {0}(-147,292)(-147,214){1}
wire w78;    //: /sn:0 {0}(-249,292)(-249,180){1}
wire w47;    //: /sn:0 {0}(441,292)(441,214){1}
wire w83;    //: /sn:0 {0}(397,534)(397,547)(365,547){1}
wire w38;    //: /sn:0 {0}(731,292)(731,222)(730,222)(730,214){1}
wire w55;    //: /sn:0 {0}(204,478)(204,439)(347,439)(347,339){1}
wire w87;    //: /sn:0 {0}(62,550)(111,550){1}
wire w43;    //: /sn:0 {0}(478,448)(478,375)(638,375)(638,339){1}
wire w9;    //: /sn:0 {0}(625,404)(673,404)(673,405)(721,405){1}
wire w79;    //: /sn:0 {0}(147,523)(147,505)(168,505){1}
wire w40;    //: /sn:0 {0}(421,504)(470,504)(470,501){1}
wire w51;    //: /sn:0 {0}(485,292)(485,180){1}
wire w57;    //: /sn:0 {0}(264,292)(264,180){1}
wire w77;    //: /sn:0 {0}(-220,292)(-220,222)(-221,222)(-221,214){1}
//: enddecls

  assign w71 = B[3]; //: TAP g44 @(-73,208) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  assign w34 = A[1]; //: TAP g8 @(775,174) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  mAND g4 (.a(w32), .b(w27), .out0(w33));   //: @(828, 293) /sz:(68, 45) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  FA g3 (.a(w16), .b(w52), .cin(w9), .cout(w19), .S(w20));   //: @(574, 382) /sz:(50, 51) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<1 ]
  assign w69 = A[0]; //: TAP g47 @(-29,174) /sn:0 /R:1 /w:[ 1 26 25 ] /ss:1
  mAND g16 (.a(w41), .b(w11), .out0(w43));   //: @(609, 293) /sz:(68, 45) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  mAND g17 (.a(w44), .b(w45), .out0(w46));   //: @(537, 293) /sz:(68, 45) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  mAND g26 (.a(w65), .b(w66), .out0(w67));   //: @(24, 293) /sz:(68, 45) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  HA g2 (.N(w46), .cin(w37), .cout(w9), .S(w21));   //: @(722, 382) /sz:(58, 49) /sn:0 /p:[ Ti0>0 Ri0>0 Lo0<1 Bo0<1 ]
  mAND g23 (.a(w59), .b(w60), .out0(w13));   //: @(171, 293) /sz:(68, 45) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  mAND g30 (.a(w74), .b(w75), .out0(w8));   //: @(-196, 293) /sz:(68, 45) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  assign w57 = A[0]; //: TAP g39 @(264,174) /sn:0 /R:1 /w:[ 1 18 17 ] /ss:1
  assign w45 = A[0]; //: TAP g24 @(556,174) /sn:0 /R:1 /w:[ 1 10 9 ] /ss:1
  //: IN g1 (B) @(-291,210) /sn:0 /w:[ 0 ]
  assign w59 = B[2]; //: TAP g60 @(220,208) /sn:0 /R:1 /w:[ 1 13 14 ] /ss:1
  assign out = {w80, w42, w39, w31, w30, w82, w21, w33}; //: CONCAT g51  @(241,667) /sn:0 /R:3 /w:[ 1 1 1 1 1 0 0 0 0 ] /dr:1 /tp:0 /drp:1
  assign w50 = B[1]; //: TAP g18 @(514,208) /sn:0 /R:1 /w:[ 1 21 22 ] /ss:1
  assign w54 = A[3]; //: TAP g10 @(338,174) /sn:0 /R:1 /w:[ 1 16 15 ] /ss:1
  mAND g25 (.a(w62), .b(w63), .out0(w12));   //: @(97, 293) /sz:(68, 45) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  assign w75 = A[2]; //: TAP g49 @(-176,174) /sn:0 /R:1 /w:[ 1 30 29 ] /ss:1
  HA g6 (.N(w7), .cin(w24), .cout(w80), .S(w42));   //: @(-109, 530) /sz:(58, 49) /sn:0 /p:[ Ti0>0 Ri0>0 Lo0<0 Bo0<0 ]
  assign w78 = A[3]; //: TAP g50 @(-249,174) /sn:0 /R:1 /w:[ 1 32 31 ] /ss:1
  FA g56 (.a(w49), .b(w70), .cin(w83), .cout(w17), .S(w30));   //: @(314, 525) /sz:(50, 51) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<1 ]
  assign w62 = B[2]; //: TAP g58 @(146,208) /sn:0 /R:1 /w:[ 1 11 12 ] /ss:1
  assign w51 = A[1]; //: TAP g9 @(485,174) /sn:0 /R:1 /w:[ 1 12 11 ] /ss:1
  assign w11 = A[3]; //: TAP g35 @(629,174) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  assign w27 = A[0]; //: TAP g7 @(848,174) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  FA g59 (.a(w79), .b(w10), .cin(w84), .cout(w87), .S(w31));   //: @(112, 524) /sz:(50, 51) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  mAND g22 (.a(w56), .b(w57), .out0(w58));   //: @(244, 293) /sz:(68, 45) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  mAND g31 (.a(w77), .b(w78), .out0(w7));   //: @(-269, 293) /sz:(68, 45) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  FA g54 (.a(w43), .b(w14), .cin(w22), .cout(w29), .S(w40));   //: @(443, 449) /sz:(50, 51) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<1 ]
  assign w74 = B[3]; //: TAP g45 @(-147,208) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  assign w63 = A[2]; //: TAP g41 @(117,174) /sn:0 /R:1 /w:[ 1 22 21 ] /ss:1
  assign w47 = B[1]; //: TAP g36 @(441,208) /sn:0 /R:1 /w:[ 1 19 20 ] /ss:1
  assign w41 = B[0]; //: TAP g33 @(657,208) /sn:0 /R:1 /w:[ 1 25 26 ] /ss:1
  FA g52 (.a(w19), .b(w58), .cin(w20), .cout(w22), .S(w82));   //: @(528, 447) /sz:(50, 51) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>0 Lo0<1 Bo0<1 ]
  assign w66 = A[3]; //: TAP g42 @(44,174) /sn:0 /R:1 /w:[ 1 24 23 ] /ss:1
  assign w60 = A[1]; //: TAP g40 @(191,174) /sn:0 /R:1 /w:[ 1 20 19 ] /ss:1
  mAND g12 (.a(w35), .b(w34), .out0(w37));   //: @(755, 293) /sz:(68, 45) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  FA g57 (.a(w55), .b(w12), .cin(w17), .cout(w79), .S(w84));   //: @(169, 479) /sz:(50, 51) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  assign w77 = B[3]; //: TAP g46 @(-221,208) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  assign w2 = A[2]; //: TAP g34 @(702,174) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  mAND g28 (.a(w71), .b(w72), .out0(w10));   //: @(-122, 293) /sz:(68, 45) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  assign w65 = B[2]; //: TAP g11 @(73,208) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:1
  assign w32 = B[0]; //: TAP g5 @(877,213) /sn:0 /R:3 /w:[ 1 32 31 ] /ss:0
  mAND g14 (.a(w38), .b(w2), .out0(w16));   //: @(682, 293) /sz:(68, 45) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  assign w56 = B[2]; //: TAP g61 @(293,208) /sn:0 /R:1 /w:[ 1 15 16 ] /ss:1
  mAND g19 (.a(w47), .b(w48), .out0(w14));   //: @(392, 293) /sz:(68, 45) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  mAND g21 (.a(w53), .b(w54), .out0(w55));   //: @(318, 293) /sz:(68, 45) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  assign w38 = B[0]; //: TAP g32 @(730,208) /sn:0 /R:1 /w:[ 1 27 28 ] /ss:1
  mAND g20 (.a(w50), .b(w51), .out0(w52));   //: @(465, 293) /sz:(68, 45) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  FA g63 (.a(w67), .b(w8), .cin(w87), .cout(w24), .S(w39));   //: @(11, 528) /sz:(50, 51) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  assign w68 = B[3]; //: TAP g43 @(-1,208) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  assign w44 = B[1]; //: TAP g15 @(586,208) /sn:0 /R:1 /w:[ 1 23 24 ] /ss:1
  //: IN g0 (A) @(-291,176) /sn:0 /w:[ 33 ]
  //: OUT g38 (out) @(298,689) /sn:0 /w:[ 0 ]
  assign w72 = A[1]; //: TAP g48 @(-102,174) /sn:0 /R:1 /w:[ 1 28 27 ] /ss:1
  mAND g27 (.a(w68), .b(w69), .out0(w70));   //: @(-49, 293) /sz:(68, 45) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  assign w53 = B[1]; //: TAP g62 @(366,208) /sn:0 /R:1 /w:[ 1 17 18 ] /ss:1
  assign w48 = A[2]; //: TAP g37 @(411,174) /sn:0 /R:1 /w:[ 1 14 13 ] /ss:1
  FA g55 (.a(w29), .b(w13), .cin(w40), .cout(w49), .S(w83));   //: @(370, 482) /sz:(50, 51) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  assign w35 = B[0]; //: TAP g13 @(803,208) /sn:0 /R:1 /w:[ 1 29 30 ] /ss:1

endmodule
//: /netlistEnd

